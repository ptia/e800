module hello;
    initial
        $display("hello, world!");
endmodule
